module mux ();
    
endmodule